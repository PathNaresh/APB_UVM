
`include "uvm_macros.svh"
import uvm_pkg::*;

`include "tb/apb_top.sv"
`include "rtl/apb_design.sv"
`include "tb/apb_intf.sv"
`include "tb/apb_pkg.sv"
