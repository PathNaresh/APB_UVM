
`include "apb_cfg.sv"
`include "apb_seq_item.sv"
`include "apb_sequence.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_scoreboard.sv"
`include "apb_agent.sv"
`include "apb_env.sv"
`include "apb_test.sv"
